/* INSERT NAME AND PENNKEY HERE */

`timescale 1ns / 1ps

`default_nettype none

/*
module lc4_alu_ctl(input  wire [15:0] i_insn
                  output wire [5:0] alu_ctl);
      // TODO
      alu_ctl[]


end module;
*/


module lc4_alu(input  wire [15:0] i_insn,
               input wire [15:0]  i_pc,
               input wire [15:0]  i_r1data,
               input wire [15:0]  i_r2data,
               output wire [15:0] o_result);


      /*** YOUR CODE HERE ***/

endmodule
